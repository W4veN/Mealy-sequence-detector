-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- Created on Wed Jan 06 09:01:23 2021

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY detector IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        R : OUT STD_LOGIC
    );
END detector;

ARCHITECTURE BEHAVIOR OF detector IS
    TYPE type_fstate IS (A,B,C,D,E,F,G);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_R : STD_LOGIC := '0';
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x,reg_R)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= A;
            reg_R <= '0';
            R <= '0';
        ELSE
            reg_R <= '0';
            R <= '0';
            CASE fstate IS
                WHEN A =>
                    IF ((x = '1')) THEN
                        reg_fstate <= B;
                    ELSIF (NOT((x = '1'))) THEN
                        reg_fstate <= C;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= A;
                    END IF;
                WHEN B =>
                    IF (NOT((x = '1'))) THEN
                        reg_fstate <= D;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= B;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= B;
                    END IF;
                WHEN C =>
                    IF ((x = '1')) THEN
                        reg_fstate <= E;
                    ELSIF (NOT((x = '1'))) THEN
                        reg_fstate <= C;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= C;
                    END IF;
                WHEN D =>
                    IF (NOT((x = '1'))) THEN
                        reg_fstate <= C;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= G;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= D;
                    END IF;
                WHEN E =>
                    IF (NOT((x = '1'))) THEN
                        reg_fstate <= F;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= B;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E;
                    END IF;
                WHEN F =>
                    IF (NOT((x = '1'))) THEN
                        reg_fstate <= C;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= G;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= F;
                    END IF;

                    IF ((x = '1')) THEN
                        reg_R <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_R <= '0';
                    END IF;
                WHEN G =>
                    IF (NOT((x = '1'))) THEN
                        reg_fstate <= F;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= B;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= G;
                    END IF;

                    IF ((x = '1')) THEN
                        reg_R <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_R <= '0';
                    END IF;
                WHEN OTHERS => 
                    reg_R <= 'X';
                    report "Reach undefined state";
            END CASE;
            R <= reg_R;
        END IF;
    END PROCESS;
END BEHAVIOR;
